/*
	Author: Quyet Luu
	Date: 7/26/2016
*/

module lab1_part6(SW,LEDR,HEX7,HEX6,HEX5,HEX4,HEX3,HEX2,HEX1,HEX0);
input [9:7] SW;
output [9:7] LEDR;
output [6:0] HEX7,HEX6,HEX5,HEX4,HEX3,HEX2,HEX1,HEX0;
reg [55:0] hex;

assign {HEX7,HEX6,HEX5,HEX4,HEX3,HEX2,HEX1,HEX0} = hex[55:0];


assign LEDR = SW; // show value of SW

always @(SW)
begin
	case(SW[9:7])
		3'h0: hex = (55'b0100001_0000110_0100100) |  ~55'b1111111_1111111_1111111;
		3'h1: hex = (55'b0100001_0000110_0100100 << 7) |  ~(55'b1111111_1111111_1111111 << 7);
		3'h2: hex = (55'b0100001_0000110_0100100 << 14) |  ~(55'b1111111_1111111_1111111 << 14);
		3'h3: hex = (55'b0100001_0000110_0100100 << 21) |  ~(55'b1111111_1111111_1111111 << 21);
		3'h4: hex = (55'b0100001_0000110_0100100 << 28) |  ~(55'b1111111_1111111_1111111 << 28);
		3'h5: hex = (55'b0100001_0000110_0100100 << 35) |  ~(55'b1111111_1111111_1111111 << 35);
		3'h6: hex = (55'b0100001_0000110_0100100 << 42 | 55'b0100001_0000110_0100100 >> 14) |  ~(55'b1111111_1111111_1111111 << 42 | 55'b1111111_1111111_1111111 >> 14 ) ;
		3'h7: hex = (55'b0100001_0000110_0100100 << 49 | 55'b0100001_0000110_0100100 >> 7) |  ~(55'b1111111_1111111_1111111 << 49 | 55'b1111111_1111111_1111111 >> 7);
		default: hex = ~(42'b0);
	endcase
end


endmodule